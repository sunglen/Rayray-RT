import(<kernel.cdl>);

celltype tInitializeRoutineBody{
	entry sRoutineBody eInitializeRoutineBody;
	call  sRoutineBody cInitialize[]; 
};
